module ansi
